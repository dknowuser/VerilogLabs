library verilog;
use verilog.vl_types.all;
entity lab1v is
end lab1v;
